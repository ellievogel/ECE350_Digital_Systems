// Author: Ellie Vogel (eov2)

module and_32();

endmodule