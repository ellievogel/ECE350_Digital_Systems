// Author: Ellie Vogel (eov2)

module and_32_bits(result, A, B);

    input [7:0] A, B;
    output [7:0] result;

    and and_gate0(result[0], A[0], B[0]);
    and and_gate1(result[1], A[1], B[1]);
    and and_gate2(result[2], A[2], B[2]);
    and and_gate3(result[3], A[3], B[3]);
    and and_gate4(result[4], A[4], B[4]);
    and and_gate5(result[5], A[5], B[5]);
    and and_gate6(result[6], A[6], B[6]);
    and and_gate7(result[7], A[7], B[7]);
    // and and_gate8(result[8], A[8], B[8]);
    // and and_gate9(result[9], A[9], B[9]);
    // and and_gate10(result[10], A[10], B[10]);
    // and and_gate11(result[11], A[11], B[11]);
    // and and_gate12(result[12], A[12], B[12]);
    // and and_gate13(result[13], A[13], B[13]);
    // and and_gate14(result[14], A[14], B[14]);
    // and and_gate15(result[15], A[15], B[15]);
    // and and_gate16(result[16], A[16], B[16]);
    // and and_gate17(result[17], A[17], B[17]);
    // and and_gate18(result[18], A[18], B[18]);
    // and and_gate19(result[19], A[19], B[19]);
    // and and_gate20(result[20], A[20], B[20]);
    // and and_gate21(result[21], A[21], B[21]);
    // and and_gate22(result[22], A[22], B[22]);
    // and and_gate23(result[23], A[23], B[23]);
    // and and_gate24(result[24], A[24], B[24]);
    // and and_gate25(result[25], A[25], B[25]);
    // and and_gate26(result[26], A[26], B[26]);
    // and and_gate27(result[27], A[27], B[27]);
    // and and_gate28(result[28], A[28], B[28]);
    // and and_gate29(result[29], A[29], B[29]);
    // and and_gate30(result[30], A[30], B[30]);
    // and and_gate31(result[31], A[31], B[31]);
endmodule