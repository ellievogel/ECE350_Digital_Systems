// Author: Ellie Vogel (eov2)

module or_32();

endmodule